/*
 * AlphaAHB V5 CPU Softcore - Advanced Vector and AI/ML Units
 * 
 * This file contains the sophisticated vector processing and AI/ML
 * acceleration units that embrace the full complexity of the
 * AlphaAHB V5 architecture.
 */

package alphaahb_v5_vector_pkg;

    // ============================================================================
    // Vector Data Types
    // ============================================================================
    
    // Explicit packed vectors for synthesis compatibility (matching Core ports)
    typedef logic [511:0] vector_512_t;  // 512-bit vector (8x64-bit FP64 elements)
    typedef logic [511:0] ai_vector_t;   // AI/ML vector (16x32-bit FP32 elements)

endpackage

// ============================================================================
// Advanced Vector Processing Unit with 512-bit SIMD (FP64)
// ============================================================================

module AdvancedVectorUnit (
    input  alphaahb_v5_vector_pkg::vector_512_t v1_data,
    input  alphaahb_v5_vector_pkg::vector_512_t v2_data,
    input  logic [3:0]  funct,
    input  logic [7:0]  mask,  // Element mask
    output alphaahb_v5_vector_pkg::vector_512_t result,
    output logic        valid,
    output logic        exception
);

    // Internal signals
    alphaahb_v5_vector_pkg::vector_512_t temp_result;
    real sum_real;
    logic valid_op;
    logic exc_flag;
    
    always_comb begin
        temp_result = 512'h0;
        valid_op = 1'b0;
        exc_flag = 1'b0;
        sum_real = 0.0;
        
        case (funct)
            4'h0: begin // VADD - Vector Addition (FP64)
                for (int i = 0; i < 8; i++) begin
                    if (mask[i]) begin
                        real r1 = $bitstoreal(v1_data[i*64 +: 64]);
                        real r2 = $bitstoreal(v2_data[i*64 +: 64]);
                        temp_result[i*64 +: 64] = $realtobits(r1 + r2);
                    end else begin
                        temp_result[i*64 +: 64] = v1_data[i*64 +: 64];
                    end
                end
                valid_op = 1'b1;
            end
            4'h1: begin // VSUB - Vector Subtraction (FP64)
                for (int i = 0; i < 8; i++) begin
                    if (mask[i]) begin
                        real r1 = $bitstoreal(v1_data[i*64 +: 64]);
                        real r2 = $bitstoreal(v2_data[i*64 +: 64]);
                        temp_result[i*64 +: 64] = $realtobits(r1 - r2);
                    end else begin
                        temp_result[i*64 +: 64] = v1_data[i*64 +: 64];
                    end
                end
                valid_op = 1'b1;
            end
            4'h2: begin // VMUL - Vector Multiplication (FP64)
                for (int i = 0; i < 8; i++) begin
                    if (mask[i]) begin
                        real r1 = $bitstoreal(v1_data[i*64 +: 64]);
                        real r2 = $bitstoreal(v2_data[i*64 +: 64]);
                        temp_result[i*64 +: 64] = $realtobits(r1 * r2);
                    end else begin
                        temp_result[i*64 +: 64] = v1_data[i*64 +: 64];
                    end
                end
                valid_op = 1'b1;
            end
            4'h3: begin // VDIV - Vector Division (FP64)
                for (int i = 0; i < 8; i++) begin
                    real r1 = $bitstoreal(v1_data[i*64 +: 64]);
                    real r2 = $bitstoreal(v2_data[i*64 +: 64]);
                    if (mask[i] && r2 != 0.0) begin
                        temp_result[i*64 +: 64] = $realtobits(r1 / r2);
                    end else begin
                        temp_result[i*64 +: 64] = v1_data[i*64 +: 64];
                    end
                end
                valid_op = 1'b1;
            end
            4'h4: begin // VFMA - Vector Fused Multiply-Add (FP64)
                for (int i = 0; i < 8; i++) begin
                    if (mask[i]) begin
                        real r1 = $bitstoreal(v1_data[i*64 +: 64]);
                        real r2 = $bitstoreal(v2_data[i*64 +: 64]);
                        // Accumulate on top of r1 (destination)
                        temp_result[i*64 +: 64] = $realtobits(r1 * r2 + r1);
                    end else begin
                        temp_result[i*64 +: 64] = v1_data[i*64 +: 64];
                    end
                end
                valid_op = 1'b1;
            end
            4'h5: begin // VREDUCE - Vector Reduction (Sum FP64)
                sum_real = 0.0;
                for (int i = 0; i < 8; i++) begin
                    real r = $bitstoreal(v1_data[i*64 +: 64]);
                    sum_real += r;
                end
                for (int i = 0; i < 8; i++) begin
                    temp_result[i*64 +: 64] = $realtobits(sum_real);
                end
                valid_op = 1'b1;
            end
            4'h6: begin // VGATHER
                for (int i = 0; i < 8; i++) begin
                    logic [2:0] idx = v2_data[i*64 +: 3];
                    if (mask[i]) begin
                        temp_result[i*64 +: 64] = v1_data[{idx, 6'b0} +: 64];
                    end else begin
                        temp_result[i*64 +: 64] = v1_data[i*64 +: 64];
                    end
                end
                valid_op = 1'b1;
            end
            4'h7: begin // VSCATTER
                temp_result = 512'h0;
                for (int i = 0; i < 8; i++) begin
                    if (mask[i]) begin
                        logic [2:0] dst_idx = v2_data[i*64 +: 3];
                        temp_result[{dst_idx, 6'b0} +: 64] = v1_data[i*64 +: 64];
                    end
                end
                valid_op = 1'b1;
            end
            4'h8: begin // VSHUFFLE
                for (int i = 0; i < 8; i++) begin
                    logic [2:0] idx = v2_data[i*64 +: 3];
                    temp_result[i*64 +: 64] = v1_data[{idx, 6'b0} +: 64];
                end
                valid_op = 1'b1;
            end
            4'h9: begin // VPERMUTE
                for (int i = 0; i < 8; i++) begin
                    logic [2:0] idx = v2_data[i*64 +: 3];
                    temp_result[i*64 +: 64] = v1_data[{idx, 6'b0} +: 64];
                end
                valid_op = 1'b1;
            end
            4'hA: begin // VBLEND
                for (int i = 0; i < 8; i++) begin
                    temp_result[i*64 +: 64] = mask[i] ? v1_data[i*64 +: 64] : v2_data[i*64 +: 64];
                end
                valid_op = 1'b1;
            end
            4'hB: begin // VSHIFT (Integer shift on 64-bit word)
                for (int i = 0; i < 8; i++) begin
                    temp_result[i*64 +: 64] = v1_data[i*64 +: 64] << v2_data[i*64 +: 6];
                end
                valid_op = 1'b1;
            end
            4'hC: begin // VROTATE (Integer rotate)
                for (int i = 0; i < 8; i++) begin
                     logic [63:0] val = v1_data[i*64 +: 64];
                     logic [5:0] rot = v2_data[i*64 +: 6];
                     temp_result[i*64 +: 64] = (val << rot) | (val >> (64 - rot));
                end
                valid_op = 1'b1;
            end
            4'hD: begin // VCOMPRESS
                int j = 0;
                for (int i = 0; i < 8; i++) begin
                    if (mask[i]) begin
                        temp_result[j*64 +: 64] = v1_data[i*64 +: 64];
                        j++;
                    end
                end
                valid_op = 1'b1;
            end
            4'hE: begin // VEXPAND
                int j = 0;
                for (int i = 0; i < 8; i++) begin
                    if (mask[i]) begin
                        temp_result[i*64 +: 64] = v1_data[j*64 +: 64];
                        j++;
                    end else begin
                        temp_result[i*64 +: 64] = 64'h0;
                    end
                end
                valid_op = 1'b1;
            end
            4'hF: begin // VCONV
                for (int i = 0; i < 8; i++) begin
                    if (mask[i]) begin
                        case (v2_data[i*64 +: 4])
                            4'h0: begin // I64->F64
                                real r = real'($signed(v1_data[i*64 +: 64]));
                                temp_result[i*64 +: 64] = $realtobits(r);
                            end
                            4'h1: begin // F64->I64
                                real r = $bitstoreal(v1_data[i*64 +: 64]);
                                temp_result[i*64 +: 64] = longint'(r);
                            end
                            4'h2: begin // F32->F64
                                real r = $bitstoshortreal(v1_data[i*64 +: 32]);
                                temp_result[i*64 +: 64] = $realtobits(r);
                            end
                            4'h3: begin // U64->F64
                                real r = real'(v1_data[i*64 +: 64]);
                                temp_result[i*64 +: 64] = $realtobits(r);
                            end
                            default: temp_result[i*64 +: 64] = v1_data[i*64 +: 64];
                        endcase
                    end else begin
                         temp_result[i*64 +: 64] = v1_data[i*64 +: 64];
                    end
                end
                valid_op = 1'b1;
            end
            default: valid_op = 1'b0;
        endcase
    end
    
    assign result = temp_result;
    assign valid = valid_op;
    assign exception = exc_flag;

endmodule

// ============================================================================
// Advanced AI/ML Unit with Neural Network Acceleration (FP32)
// ============================================================================

module AdvancedAIMLUnit (
    input  logic        clk,
    input  logic        rst_n,
    input  alphaahb_v5_vector_pkg::ai_vector_t input_data,
    input  alphaahb_v5_vector_pkg::ai_vector_t weight_data,
    input  alphaahb_v5_vector_pkg::ai_vector_t bias_data,
    input  alphaahb_v5_vector_pkg::vector_512_t state_data, // Added for stateful ops
    input  logic [3:0]  funct,
    input  logic [7:0]  config,
    output alphaahb_v5_vector_pkg::ai_vector_t result,
    output logic        valid,
    output logic        exception
);

    alphaahb_v5_vector_pkg::ai_vector_t temp_result;
    real sum_accum;
    real exp_val_buf [15:0];
    real sum_exp;
    logic valid_op;
    logic exc_flag;

    // Stateful LFSR for Dropout
    logic [15:0] lfsr_reg;
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            lfsr_reg <= 16'hACE1;
        end else begin
            // Free-running LFSR (Galois or Fibonacci)
            // Taps: 16, 14, 13, 11 (Xilinx xapp) -> indices 15, 13, 12, 10
            logic feedback = lfsr_reg[15] ^ lfsr_reg[13] ^ lfsr_reg[12] ^ lfsr_reg[10];
            lfsr_reg <= {lfsr_reg[14:0], feedback};
        end
    end
    
    always_comb begin
        temp_result = 512'h0;
        valid_op = 1'b0;
        exc_flag = 1'b0;
        sum_accum = 0.0;
        sum_exp = 0.0;
        
        case (funct)
            4'h0: begin // CONV - Convolution Operation (FP32)
                for (int i = 0; i < 16; i++) begin
                    sum_accum = 0.0;
                    for (int j = 0; j < 16; j++) begin
                        shortreal i_val = $bitstoshortreal(input_data[j*32 +: 32]);
                        shortreal w_val = $bitstoshortreal(weight_data[j*32 +: 32]);
                        sum_accum += (i_val * w_val);
                    end
                    // Add bias
                    shortreal b_val = $bitstoshortreal(bias_data[i*32 +: 32]);
                    temp_result[i*32 +: 32] = $shortrealtobits(shortreal'(sum_accum) + b_val);
                end
                valid_op = 1'b1;
            end
            4'h1: begin // FC - Fully Connected (FP32)
                for (int i = 0; i < 16; i++) begin
                    sum_accum = 0.0;
                    for (int j = 0; j < 16; j++) begin
                        shortreal i_val = $bitstoshortreal(input_data[j*32 +: 32]);
                        shortreal w_val = $bitstoshortreal(weight_data[j*32 +: 32]);
                        sum_accum += (i_val * w_val);
                    end
                    shortreal b_val = $bitstoshortreal(bias_data[i*32 +: 32]);
                    temp_result[i*32 +: 32] = $shortrealtobits(shortreal'(sum_accum) + b_val);
                end
                valid_op = 1'b1;
            end
            4'h2: begin // RELU (FP32)
                for (int i = 0; i < 16; i++) begin
                    shortreal val = $bitstoshortreal(input_data[i*32 +: 32]);
                    temp_result[i*32 +: 32] = (val > 0.0) ? input_data[i*32 +: 32] : 32'h0;
                end
                valid_op = 1'b1;
            end
            4'h3: begin // SIGMOID (FP32 Pade)
                for (int i = 0; i < 16; i++) begin
                    real x_val = $bitstoshortreal(input_data[i*32 +: 32]);
                    real sigmoid_result;
                    if (x_val >= 10.0) sigmoid_result = 1.0;
                    else if (x_val <= -10.0) sigmoid_result = 0.0;
                    else begin
                        real x2 = x_val * x_val;
                        real x4 = x2 * x2;
                        real P = 0.5 + 0.25 * x2 + 0.0125 * x4;
                        real Q = 1.0 + 1.0 * x2 + 0.25 * x4;
                        sigmoid_result = 0.5 + x_val * (P / Q);
                    end
                    temp_result[i*32 +: 32] = $shortrealtobits(shortreal'(sigmoid_result));
                end
                valid_op = 1'b1;
            end
            4'h4: begin // TANH
                for (int i = 0; i < 16; i++) begin
                    real x_val = $bitstoshortreal(input_data[i*32 +: 32]);
                    real x2 = 2.0 * x_val;
                    real sig2;
                    if (x2 >= 10.0) sig2 = 1.0;
                    else if (x2 <= -10.0) sig2 = 0.0;
                    else begin
                        real x2sq = x2 * x2;
                        real x4sq = x2sq * x2sq;
                        real P = 0.5 + 0.25 * x2sq + 0.0125 * x4sq;
                        real Q = 1.0 + 1.0 * x2sq + 0.25 * x4sq;
                        sig2 = 0.5 + x2 * (P / Q);
                    end
                    temp_result[i*32 +: 32] = $shortrealtobits(shortreal'(2.0 * sig2 - 1.0));
                end
                valid_op = 1'b1;
            end
            4'h5: begin // SOFTMAX
                shortreal max_val = $bitstoshortreal(input_data[0 +: 32]);
                for (int i = 1; i < 16; i++) begin
                    shortreal val = $bitstoshortreal(input_data[i*32 +: 32]);
                    if (val > max_val) max_val = val;
                end
                
                sum_exp = 0.0;
                for (int i = 0; i < 16; i++) begin
                    real x_val = $bitstoshortreal(input_data[i*32 +: 32]);
                    real shifted = x_val - max_val;
                    if (shifted > 10.0) shifted = 10.0;
                    else if (shifted < -10.0) shifted = -10.0;
                    exp_val_buf[i] = $exp(shifted);
                    sum_exp += exp_val_buf[i];
                end
                
                for (int i = 0; i < 16; i++) begin
                    temp_result[i*32 +: 32] = $shortrealtobits(shortreal'(exp_val_buf[i] / sum_exp));
                end
                valid_op = 1'b1;
            end
            4'h6: begin // POOL
                int pool_size = (config[3:0] == 0) ? 2 : config[3:0];
                int pool_type = config[7:4];
                
                for (int i = 0; i < 16; i += pool_size) begin
                    real p_res = $bitstoshortreal(input_data[i*32 +: 32]);
                    int count = 1;
                    
                    for (int j = 1; j < pool_size && (i+j) < 16; j++) begin
                        real c = $bitstoshortreal(input_data[(i+j)*32 +: 32]);
                        count++;
                        if (pool_type == 0) begin if (c > p_res) p_res = c; end // Max
                        else if (pool_type == 1) p_res += c; // Avg (step 1)
                        else if (pool_type == 2) begin if (c < p_res) p_res = c; end // Min
                    end
                    
                    if (pool_type == 1) p_res = p_res / count;
                    
                    for (int j = 0; j < pool_size && (i+j) < 16; j++) begin
                        temp_result[(i+j)*32 +: 32] = $shortrealtobits(shortreal'(p_res));
                    end
                end
                valid_op = 1'b1;
            end
            4'h7: begin // BATCHNORM
                // Calculate Mean
                sum_accum = 0.0;
                for (int i = 0; i < 16; i++) sum_accum += $bitstoshortreal(input_data[i*32 +: 32]);
                real mean_val = sum_accum / 16.0;
                
                // Calculate Variance (2nd pass)
                real var_accum = 0.0;
                for (int i = 0; i < 16; i++) begin
                    real val = $bitstoshortreal(input_data[i*32 +: 32]);
                    real diff = val - mean_val;
                    var_accum += diff * diff;
                end
                real variance = var_accum / 16.0;
                // Calculate Inverse Stdev with Epsilon
                real inv_std = 1.0 / $sqrt(variance + 1.0e-5); 
                
                for (int i = 0; i < 16; i++) begin
                    real val = $bitstoshortreal(input_data[i*32 +: 32]);
                    real norm = (val - mean_val) * inv_std;
                    real w = $bitstoshortreal(weight_data[i*32 +: 32]);
                    real b = $bitstoshortreal(bias_data[i*32 +: 32]);
                    temp_result[i*32 +: 32] = $shortrealtobits(shortreal'(norm * w + b));
                end
                valid_op = 1'b1;
            end
            4'h8: begin // DROPOUT
                // Use stateful LFSR
                logic [15:0] lfsr_temp = lfsr_reg;
                logic [7:0] keep_prob = config;
                real scale = 256.0 / (real'(keep_prob) + 1.0);
                
                for (int i = 0; i < 16; i++) begin
                    // Compute pseudo-random value for this element
                    logic feedback = lfsr_temp[15] ^ lfsr_temp[13] ^ lfsr_temp[12] ^ lfsr_temp[10];
                    lfsr_temp = {lfsr_temp[14:0], feedback};
                    
                    logic [7:0] rand_val = lfsr_temp[7:0]; 
                    if (rand_val < keep_prob) begin
                         real val = $bitstoshortreal(input_data[i*32 +: 32]);
                         temp_result[i*32 +: 32] = $shortrealtobits(shortreal'(val * scale));
                    end else begin
                         temp_result[i*32 +: 32] = 32'h0;
                    end
                end
                valid_op = 1'b1;
            end
            4'h9: begin // LSTM (Real State)
                // Use state_data for h_{t-1}. c_{t-1} assumed 0 for instruction step context
                for (int i = 0; i < 16; i++) begin
                    real x = $bitstoshortreal(input_data[i*32 +: 32]);
                    real w = $bitstoshortreal(weight_data[i*32 +: 32]);
                    real b = $bitstoshortreal(bias_data[i*32 +: 32]);
                    real h_prev = $bitstoshortreal(state_data[i*32 +: 32]); // Use 512-bit state if available, mapping 1:1 with vector
                    
                    real pre = w * x + b + h_prev * 0.1; // Added recurrent weight equivalent
                    
                    // Gates (Same Pade logic for brevity, reused across Update/Reset/Out)
                    real sig;
                    if (pre > 10) sig = 1; else if (pre < -10) sig = 0;
                    else sig = 1.0 / (1.0 + $exp(-pre)); // Using $exp for cleanliness
                    
                    real f_g = sig; 
                    real i_g = sig; 
                    real o_g = sig;
                    real c_cand = (2.0 / (1.0 + $exp(-2.0*pre))) - 1.0; // Tanh
                    
                    real c_t = f_g * 0.0 + i_g * c_cand; // c_prev=0
                    real h_t = o_g * ((2.0 / (1.0 + $exp(-2.0*c_t))) - 1.0);
                    
                    temp_result[i*32 +: 32] = $shortrealtobits(shortreal'(h_t));
                end
                valid_op = 1'b1;
            end
            4'hA: begin // GRU (Real State)
                for (int i = 0; i < 16; i++) begin
                    real x = $bitstoshortreal(input_data[i*32 +: 32]);
                    real w = $bitstoshortreal(weight_data[i*32 +: 32]);
                    real b = $bitstoshortreal(bias_data[i*32 +: 32]);
                    real h_prev = $bitstoshortreal(state_data[i*32 +: 32]);
                    
                    real pre = w * x + b + h_prev * 0.1;
                    real z = 1.0 / (1.0 + $exp(-pre));
                    real r = 1.0 / (1.0 + $exp(-pre));
                    real h_cand = (2.0 / (1.0 + $exp(-2.0 * (w*x + r*h_prev)))) - 1.0;
                    real h_t = (1.0 - z) * h_prev + z * h_cand;
                    
                    temp_result[i*32 +: 32] = $shortrealtobits(shortreal'(h_t));
                end
                valid_op = 1'b1;
            end
            4'hB: begin // ATTENTION
                 // Vector Attention: Softmax(Input * Weight) * Bias
                 // Interpreted as: Element-wise score, then normalize, then scale.
                 real scale = 0.25; // 1/sqrt(16)
                 for (int i = 0; i < 16; i++) begin
                     real q = $bitstoshortreal(input_data[i*32 +: 32]);
                     real k = $bitstoshortreal(weight_data[i*32 +: 32]);
                     exp_val_buf[i] = q * k * scale;
                 end
                 // Softmax on scores
                 sum_exp = 0.0;
                 for (int i = 0; i < 16; i++) { exp_val_buf[i] = $exp(exp_val_buf[i]); sum_exp += exp_val_buf[i]; }
                 for (int i = 0; i < 16; i++) {
                     real attn = exp_val_buf[i] / sum_exp;
                     real v = $bitstoshortreal(bias_data[i*32 +: 32]); // Value from bias vector?
                     temp_result[i*32 +: 32] = $shortrealtobits(shortreal'(attn * v));
                 }
                 valid_op = 1'b1;
            end
            default: valid_op = 1'b0;
        endcase
    end
    
    assign result = temp_result;
    assign valid = valid_op;
    assign exception = exc_flag;

endmodule
